module MemoriadeInstrucoes(address,clock,instruction);

input[31:0] address;
input clock;
output [31:0] instruction;
integer flag=0;
reg[31:0] instrmem[31:0];

always @(posedge clock) begin

	if(flag==0) 
	begin
	/*//fibonacci
	   instrmem[0]= 32'b010010_00000_00000_00000_00000000000; //nop
		instrmem[1]= 32'b001100_00000_00001_00000_00000000001; // r[1]=1
		instrmem[2]= 32'b001100_00000_00010_00000_00000000001; // r[2]=1
		instrmem[3]= 32'b001100_00000_00100_00000_00000000000; // r[4]=0
		instrmem[4]= 32'b010100_00000_00000_00011_00000000000; // input
		instrmem[5]= 32'b000011_00011_00011_00000_00000000001; // r[3]=r[3]-1
		instrmem[6]= 32'b000110_00000_00011_01010_00000000000; // slt r[10],r[0],r[3]
		instrmem[7]= 32'b001110_01010_00000_00000_00000001100; // beq 12,[r10],r[0]
		instrmem[8]= 32'b000000_00001_00100_00010_00000000000; // r[2]= r[1]+r[4]
		instrmem[9]= 32'b010110_00001_00000_00100_00000000000; //r4=r1
		instrmem[10]= 32'b010110_00010_00000_00001_00000000000; //r1=r2
		instrmem[11]= 32'b010000_00000_00000_00000_00000000101; //jump to 5
		instrmem[12]= 32'b001100_00000_00101_00000_00000001111; // r[5]=15 ldi
		instrmem[13]= 32'b010001_00101_00000_00000_00000000000; // jmpr
		instrmem[15]= 32'b001101_00000_00010_00000_00000000010; // SW
		instrmem[16]= 32'b001011_00000_00110_00000_00000000010; //lw
		instrmem[17]= 32'b010101_00110_00000_00000_00000000000; // out r[2]
		instrmem[18]= 32'b010011_00000_00000_00000_00000000000; //halt*/
		
		/*			
		/// fibonacci2
		instrmem[0]= 32'b010010_00000_00000_00000_00000000000; //nop
		instrmem[1]= 32'b000010_00000_00001_00000_00000000001; // r[1]=1 addi
		instrmem[2]= 32'b001100_00000_00010_00000_00000000001; // r[2]=1 ldi
		instrmem[3]= 32'b001100_00000_00100_00000_00000000000; // r[4]=0 //ldi
		instrmem[4]= 32'b010100_00000_00000_00011_00000000000; // input 
		instrmem[5]= 32'b000001_00011_00001_00011_00000000000; // r[3]=r[3]-r[1] //sub
		instrmem[6]= 32'b000110_00000_00011_01010_00000000000; // slt r[10],r[0],r[3] //slt
		instrmem[7]= 32'b001110_01010_00000_00000_00000001101; // beq 13,[r10],r[0] //beq
		instrmem[8]= 32'b000000_00001_00100_00010_00000000000; // r[2]= r[1]+r[4] //add
		instrmem[9]= 32'b010110_00001_00000_00100_00000000000; //r4=r1 //move
		instrmem[10]= 32'b010110_00010_00000_00001_00000000000; //r1=r2 //move
		instrmem[11]= 32'b000011_00011_00011_00000_00000000001; // r[3]=r[3]-1 //subi
		instrmem[12]= 32'b010000_00000_00000_00000_00000000110; //jump to 6 //jmp
		instrmem[13]= 32'b010001_00101_00000_00000_00000000000; // jmpr //jumptoreg
		instrmem[15]= 32'b001101_00000_00010_00000_00000000010; // SW //sw
		instrmem[16]= 32'b001011_00000_00110_00000_00000000010; //lw //lw
		instrmem[17]= 32'b000111_00000_00110_00000_00000000000; //NOT
		instrmem[18]= 32'b000111_00000_00110_00000_00000000000; //NOT
		instrmem[19]= 32'b010101_00110_00000_00000_00000000000; // out r[2] //output
		instrmem[20]= 32'b010011_00000_00000_00000_00000000000; //halt 
*/
	/*	//todas instruçoes
		instrmem[0]= 32'b010100_00000_00000_00001_00000000000; // input r[1]=1
		instrmem[1]= 32'b010100_00000_00000_00010_00000000000; // input r[2]=2
		instrmem[2]= 32'b001100_00000_00100_00000_00000001111; // r[4]=15 //ldi
		instrmem[3]= 32'b000000_00001_00010_00011_00000000000; // r[3]= r[1]+r[2] //add
		instrmem[4]= 32'b000001_00001_00010_00011_00000000000; // r[3]= r[1]-r[2] //sub
		instrmem[5]= 32'b000100_00001_00010_00011_00000000000; // r[3]= r[1]*r[2] //mult
		instrmem[6]= 32'b000101_00001_00010_00011_00000000000; // r[3]= r[1]/r[2] //div
		instrmem[7]= 32'b011000_00001_00000_00001_00001_000000; // r[1]=SHFR[r1]
		instrmem[8]= 32'b010111_00010_00000_00010_00001_000000; //r[2]=SHFL[r2]
		instrmem[9]= 32'b010110_00001_00000_00011_00000000000; //r3=r1 //move
		instrmem[10]= 32'b010110_00010_00000_00001_00000000000; //r1=r2 //move
		instrmem[11]= 32'b000011_00011_00011_00000_00000000001; // r[3]=r[3]-1 //subi
		instrmem[12]= 32'b000010_00010_00010_00000_00000000001; // r[2]=r[2]+1 //addi
		instrmem[13]= 32'b010001_00100_00000_00000_00000000000; // jmpr[15]
		instrmem[15]= 32'b010010_00000_00000_00000_00000000000; //nop
		instrmem[16]= 32'b010110_00100_00000_00011_00000000000; //r3=r4 //move
		instrmem[17]= 32'b000111_00011_00000_00011_00000000000; //NOT r3
		instrmem[18]= 32'b000111_00011_00000_00011_00000000000; //NOT r3
		instrmem[19]= 32'b001000_00011_00100_00101_00000000000; // r[5]= r3 AND r4
		instrmem[20]= 32'b001001_00011_00100_00110_00000000000; // r[6]= r3 OR r4
		instrmem[21]= 32'b001010_00011_00100_00111_00000000000; // r[7]= r3 XOR r2
		instrmem[22]= 32'b001110_00101_00011_00000_00000011001; // beq 25,[r5],r[3] //beq
		instrmem[23]= 32'b010000_00000_00000_00000_00000011100; //jump to 28 //jmp
		instrmem[25]= 32'b000110_00101_00011_01010_00000000000; // slt r[10],r[5],r[3] //slt
		instrmem[26]= 32'b001111_00101_01010_00000_00000011100; // bne 28,[r5],r[10] //beq
		instrmem[28]= 32'b001101_00000_00101_00000_00000000010; // SW r[5]
		instrmem[29]= 32'b001011_00000_01000_00000_00000000010; // LW r[8]
		instrmem[30]= 32'b010101_01010_00000_00000_00000000000; // out r[10] //output
		instrmem[31]= 32'b010011_00000_00000_00000_00000000000; //halt
		*/
		
		
		
		
		
//				calcular delta com a=2, b=4 e c=1
	/*	instrmem[0]= 32'bb010100_00000_00000_00001_00000000000; // inpu
		instrmem[2]= 32'b010100_00000_00000_00010_00000000000; // input
		instrmem[4]= 32'b010100_00000_00000_00011_00000000000; // input
		instrmem[6]= 32'b001100_00000_00100_00000_00000000100; // r[4]=4
		instrmem[7]= 32'b000100_00100_00100_00010_00000000000; // b=b^2=b*b
		instrmem[8]= 32'b000100_00100_00001_00100_00000000000; // r[4]=4*a
		instrmem[9]= 32'b000100_00100_00011_00100_00000000000; // r[4]=4*a*c
		instrmem[10]= 32'b000001_00010_00100_00100_00000000000; // r[4]=b^2-4*a*c
		instrmem[11]= 32'b010101_00100_00000_00000_00000000000; // out r[4]
		instrmem[12]= 32'b010011_00000_00000_00000_00000000000; //halt*/
		
	
	// verifica se dois triangulos tem areas iguais, caso sim sai 1, caso nao sai 2
	
		/*instrmem[0]= 32'b010010_00000_00000_00000_00000000000; //nop
		instrmem[1]= 32'b010100_00000_00000_00011_00000000000; // input base r3
	   instrmem[2]= 32'b010010_00000_00000_00000_00000000000; //nop
		instrmem[3]= 32'b010010_00000_00000_00000_00000000000; //nop
		instrmem[4]= 32'b010010_00000_00000_00000_00000000000; //nop
		instrmem[5]= 32'b010100_00000_00000_00010_00000000000; // input altura r2
		instrmem[6]= 32'b000100_00010_00011_00100_00000000000; // r[4]= base*altura //MULT  r4
		instrmem[7]= 32'b010010_00000_00000_00000_00000000000; //nop
		instrmem[8]= 32'b010010_00000_00000_00000_00000000000; //nop
		instrmem[9]= 32'b010010_00000_00000_00000_00000000000; //nop
		instrmem[10]= 32'b011000_00100_00000_00100_00001_000000; // base*altura/2 - SHFR
		instrmem[11]= 32'b010111_00100_00000_00100_00001_000000; // base*altura/2 - SHFL
		instrmem[12]= 32'b001100_00000_00101_00000_00000000010; // r[5]=2 ldi   r5
		instrmem[13]= 32'b000101_00100_00101_00100_00000_000000; // r4 = base*altura/2 - div
		instrmem[14]= 32'b010010_00000_00000_00000_00000000000; //nop
		instrmem[15]= 32'b010100_00000_00000_00001_00000000000; // input base   r1
		instrmem[16]= 32'b010010_00000_00000_00000_00000000000; //nop
		instrmem[17]= 32'b010010_00000_00000_00000_00000000000; //nop
		instrmem[18]= 32'b010100_00000_00000_00110_00000000000; //input altura  r6
		instrmem[19]= 32'b000100_00001_00110_00110_00000000000; // r[6]= base*altura //MULT  r4
		instrmem[20]= 32'b000101_00110_00101_00110_00000000000; // base*altura/2 - SHFR - base*altura/2
		instrmem[21]= 32'b001000_00100_00110_00111_00000_000000; // r4 = AND r4 r6 
		instrmem[22]= 32'b001111_00110_00100_00000_00000011010; // bne 26,[r4],r[6] //bne
		instrmem[23]= 32'b000011_00101_00101_00000_00000000001; // r[5]-1 //subi
		instrmem[24]= 32'b010101_00101_00000_00000_00000000000; // out r[5]
		instrmem[25]= 32'b010011_00000_00000_00000_00000000000; //halt
		instrmem[26]= 32'b001010_00100_00110_00100_00000000000; // r4 = xor r4 r6
		instrmem[27]= 32'b001111_00100_00110_00000_00000011110; // bne 30,[r6],r[4] //bne
		instrmem[28]= 32'b010010_00000_00000_00000_00000000000; //nop
		instrmem[29]= 32'b010010_00000_00000_00000_00000000000; //nop
		instrmem[30]= 32'b010101_00101_00000_00000_00000000000; // out r[2]
		instrmem[31]= 32'b010011_00000_00000_00000_00000000000; //halt*/
		
	///nao sei
		
		/*instrmem[2]=  32'b000000_00001_00001_00100_00000000000; // r[3]= r[1]+r[1]
		instrmem[3]=   32'b001000_00001_00100_00101_00000000000; // AND
		instrmem[4]=   32'b001001_00001_00100_00110_00000000000; // OR
		instrmem[5]=   32'b001010_00001_00100_00111_00000000000; // xOR
		instrmem[2]=  32'b001101_00001_00001_00000_00000000010; // SW
		instrmem[3]=  32'b001011_00001_00010_00000_00000000010;  //lw
		instrmem[4]=  32'b010000_00000_00000_00000_00000000110;
		instrmem[6]=  32'b010001_01001_00000_00000_00000000000;  //add
		instrmem[9]=  32'b000000_00001_00001_00100_00000000000;
		instrmem[10]=  32'b000000_00001_00001_00100_00000000000;
		instrmem[11]=  32'b010010_00000_00000_00000_00000000000;
		instrmem[12]=  32'b000000_00001_00001_00100_00000000000;
		//instrmem[13]=  32'b010011_00000_00000_00000_00000000000;
		instrmem[13]=  32'b010111_01000_00000_00101_00001000000;
		instrmem[14]=  32'b011000_01000_00000_00110_00001000000;
		instrmem[15]=  32'b010110_00001_00000_00111_00000000000;
		instrmem[16]=  32'b000000_00111_00111_01000_00000000000;
		//instrmem[6]=   32'b001011_00001_00100_01111_0000000000; // XOR
		instrmem[2] = 32'b000001_00011_00001_00011_00000000000; // r[3]= r[3]-r[1]*/
		//instrmem[3] = 32'b000110_00010_00001_00011_00000000000; // r[2]= r[3]*r[3]
		//instrmem[4] = 32'b000111_00011_00000_00100_00000000101; // r[4]= r[2]/r[3] */
		flag<=1;
	end
end

assign instruction=instrmem[address];

endmodule 